-- core.vhd

-- Generated using ACDS version 16.1 196

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity core is
	port (
		clk_clk                           : in  std_logic                     := '0';             --                        clk.clk
		freq_0_external_connection_export : in  std_logic_vector(23 downto 0) := (others => '0'); -- freq_0_external_connection.export
		freq_1_external_connection_export : in  std_logic_vector(23 downto 0) := (others => '0'); -- freq_1_external_connection.export
		freq_2_external_connection_export : in  std_logic_vector(23 downto 0) := (others => '0'); -- freq_2_external_connection.export
		freq_3_external_connection_export : in  std_logic_vector(23 downto 0) := (others => '0'); -- freq_3_external_connection.export
		freq_4_external_connection_export : in  std_logic_vector(23 downto 0) := (others => '0'); -- freq_4_external_connection.export
		freq_5_external_connection_export : in  std_logic_vector(23 downto 0) := (others => '0'); -- freq_5_external_connection.export
		freq_6_external_connection_export : in  std_logic_vector(23 downto 0) := (others => '0'); -- freq_6_external_connection.export
		freq_7_external_connection_export : in  std_logic_vector(23 downto 0) := (others => '0'); -- freq_7_external_connection.export
		hum_export                        : in  std_logic_vector(15 downto 0) := (others => '0'); --                        hum.export
		pwm_0_external_connection_export  : out std_logic_vector(6 downto 0);                     --  pwm_0_external_connection.export
		pwm_1_external_connection_export  : out std_logic_vector(6 downto 0);                     --  pwm_1_external_connection.export
		pwm_2_external_connection_export  : out std_logic_vector(6 downto 0);                     --  pwm_2_external_connection.export
		pwm_3_external_connection_export  : out std_logic_vector(6 downto 0);                     --  pwm_3_external_connection.export
		pwm_4_external_connection_export  : out std_logic_vector(6 downto 0);                     --  pwm_4_external_connection.export
		pwm_5_external_connection_export  : out std_logic_vector(6 downto 0);                     --  pwm_5_external_connection.export
		pwm_6_external_connection_export  : out std_logic_vector(6 downto 0);                     --  pwm_6_external_connection.export
		pwm_7_external_connection_export  : out std_logic_vector(6 downto 0);                     --  pwm_7_external_connection.export
		tem_export                        : in  std_logic_vector(15 downto 0) := (others => '0'); --                        tem.export
		uart_external_connection_rxd      : in  std_logic                     := '0';             --   uart_external_connection.rxd
		uart_external_connection_txd      : out std_logic                                         --                           .txd
	);
end entity core;

architecture rtl of core is
	component core_Hum is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(15 downto 0) := (others => 'X')  -- export
		);
	end component core_Hum;

	component core_freq_0 is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(23 downto 0) := (others => 'X')  -- export
		);
	end component core_freq_0;

	component core_nios2_gen2_0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(15 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(15 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component core_nios2_gen2_0;

	component core_onchip_memory2_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(11 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component core_onchip_memory2_0;

	component core_pwm_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(6 downto 0)                      -- export
		);
	end component core_pwm_0;

	component core_timer_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component core_timer_0;

	component core_uart is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			read_n        : in  std_logic                     := 'X';             -- read_n
			write_n       : in  std_logic                     := 'X';             -- write_n
			writedata     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			rxd           : in  std_logic                     := 'X';             -- export
			txd           : out std_logic;                                        -- export
			irq           : out std_logic                                         -- irq
		);
	end component core_uart;

	component core_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                  : in  std_logic                     := 'X';             -- clk
			nios2_gen2_0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			nios2_gen2_0_data_master_address               : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_data_master_waitrequest           : out std_logic;                                        -- waitrequest
			nios2_gen2_0_data_master_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_gen2_0_data_master_read                  : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_data_master_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_gen2_0_data_master_write                 : in  std_logic                     := 'X';             -- write
			nios2_gen2_0_data_master_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_gen2_0_data_master_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			nios2_gen2_0_instruction_master_address        : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_instruction_master_waitrequest    : out std_logic;                                        -- waitrequest
			nios2_gen2_0_instruction_master_read           : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_instruction_master_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			freq_0_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			freq_0_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			freq_1_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			freq_1_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			freq_2_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			freq_2_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			freq_3_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			freq_3_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			freq_4_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			freq_4_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			freq_5_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			freq_5_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			freq_6_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			freq_6_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			freq_7_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			freq_7_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Hum_s1_address                                 : out std_logic_vector(1 downto 0);                     -- address
			Hum_s1_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_gen2_0_debug_mem_slave_address           : out std_logic_vector(8 downto 0);                     -- address
			nios2_gen2_0_debug_mem_slave_write             : out std_logic;                                        -- write
			nios2_gen2_0_debug_mem_slave_read              : out std_logic;                                        -- read
			nios2_gen2_0_debug_mem_slave_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_gen2_0_debug_mem_slave_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_gen2_0_debug_mem_slave_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess       : out std_logic;                                        -- debugaccess
			onchip_memory2_0_s1_address                    : out std_logic_vector(11 downto 0);                    -- address
			onchip_memory2_0_s1_write                      : out std_logic;                                        -- write
			onchip_memory2_0_s1_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_0_s1_writedata                  : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_0_s1_byteenable                 : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_0_s1_chipselect                 : out std_logic;                                        -- chipselect
			onchip_memory2_0_s1_clken                      : out std_logic;                                        -- clken
			pwm_0_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			pwm_0_s1_write                                 : out std_logic;                                        -- write
			pwm_0_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pwm_0_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			pwm_0_s1_chipselect                            : out std_logic;                                        -- chipselect
			pwm_1_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			pwm_1_s1_write                                 : out std_logic;                                        -- write
			pwm_1_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pwm_1_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			pwm_1_s1_chipselect                            : out std_logic;                                        -- chipselect
			pwm_2_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			pwm_2_s1_write                                 : out std_logic;                                        -- write
			pwm_2_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pwm_2_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			pwm_2_s1_chipselect                            : out std_logic;                                        -- chipselect
			pwm_3_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			pwm_3_s1_write                                 : out std_logic;                                        -- write
			pwm_3_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pwm_3_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			pwm_3_s1_chipselect                            : out std_logic;                                        -- chipselect
			pwm_4_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			pwm_4_s1_write                                 : out std_logic;                                        -- write
			pwm_4_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pwm_4_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			pwm_4_s1_chipselect                            : out std_logic;                                        -- chipselect
			pwm_5_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			pwm_5_s1_write                                 : out std_logic;                                        -- write
			pwm_5_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pwm_5_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			pwm_5_s1_chipselect                            : out std_logic;                                        -- chipselect
			pwm_6_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			pwm_6_s1_write                                 : out std_logic;                                        -- write
			pwm_6_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pwm_6_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			pwm_6_s1_chipselect                            : out std_logic;                                        -- chipselect
			pwm_7_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			pwm_7_s1_write                                 : out std_logic;                                        -- write
			pwm_7_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pwm_7_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			pwm_7_s1_chipselect                            : out std_logic;                                        -- chipselect
			Tem_s1_address                                 : out std_logic_vector(1 downto 0);                     -- address
			Tem_s1_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_address                             : out std_logic_vector(2 downto 0);                     -- address
			timer_0_s1_write                               : out std_logic;                                        -- write
			timer_0_s1_readdata                            : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_writedata                           : out std_logic_vector(15 downto 0);                    -- writedata
			timer_0_s1_chipselect                          : out std_logic;                                        -- chipselect
			uart_s1_address                                : out std_logic_vector(2 downto 0);                     -- address
			uart_s1_write                                  : out std_logic;                                        -- write
			uart_s1_read                                   : out std_logic;                                        -- read
			uart_s1_readdata                               : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			uart_s1_writedata                              : out std_logic_vector(15 downto 0);                    -- writedata
			uart_s1_begintransfer                          : out std_logic;                                        -- begintransfer
			uart_s1_chipselect                             : out std_logic                                         -- chipselect
		);
	end component core_mm_interconnect_0;

	component core_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component core_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal nios2_gen2_0_debug_reset_request_reset                     : std_logic;                     -- nios2_gen2_0:debug_reset_request -> [rst_controller:reset_in0, rst_controller:reset_in1]
	signal nios2_gen2_0_data_master_readdata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	signal nios2_gen2_0_data_master_waitrequest                       : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	signal nios2_gen2_0_data_master_debugaccess                       : std_logic;                     -- nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	signal nios2_gen2_0_data_master_address                           : std_logic_vector(15 downto 0); -- nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	signal nios2_gen2_0_data_master_byteenable                        : std_logic_vector(3 downto 0);  -- nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	signal nios2_gen2_0_data_master_read                              : std_logic;                     -- nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	signal nios2_gen2_0_data_master_write                             : std_logic;                     -- nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	signal nios2_gen2_0_data_master_writedata                         : std_logic_vector(31 downto 0); -- nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	signal nios2_gen2_0_instruction_master_readdata                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	signal nios2_gen2_0_instruction_master_waitrequest                : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	signal nios2_gen2_0_instruction_master_address                    : std_logic_vector(15 downto 0); -- nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	signal nios2_gen2_0_instruction_master_read                       : std_logic;                     -- nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata    : std_logic_vector(31 downto 0); -- nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest : std_logic;                     -- nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address     : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read        : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable  : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write       : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata   : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	signal mm_interconnect_0_timer_0_s1_chipselect                    : std_logic;                     -- mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	signal mm_interconnect_0_timer_0_s1_readdata                      : std_logic_vector(15 downto 0); -- timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	signal mm_interconnect_0_timer_0_s1_address                       : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_0_s1_address -> timer_0:address
	signal mm_interconnect_0_timer_0_s1_write                         : std_logic;                     -- mm_interconnect_0:timer_0_s1_write -> mm_interconnect_0_timer_0_s1_write:in
	signal mm_interconnect_0_timer_0_s1_writedata                     : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	signal mm_interconnect_0_freq_7_s1_readdata                       : std_logic_vector(31 downto 0); -- freq_7:readdata -> mm_interconnect_0:freq_7_s1_readdata
	signal mm_interconnect_0_freq_7_s1_address                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:freq_7_s1_address -> freq_7:address
	signal mm_interconnect_0_freq_6_s1_readdata                       : std_logic_vector(31 downto 0); -- freq_6:readdata -> mm_interconnect_0:freq_6_s1_readdata
	signal mm_interconnect_0_freq_6_s1_address                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:freq_6_s1_address -> freq_6:address
	signal mm_interconnect_0_freq_5_s1_readdata                       : std_logic_vector(31 downto 0); -- freq_5:readdata -> mm_interconnect_0:freq_5_s1_readdata
	signal mm_interconnect_0_freq_5_s1_address                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:freq_5_s1_address -> freq_5:address
	signal mm_interconnect_0_freq_4_s1_readdata                       : std_logic_vector(31 downto 0); -- freq_4:readdata -> mm_interconnect_0:freq_4_s1_readdata
	signal mm_interconnect_0_freq_4_s1_address                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:freq_4_s1_address -> freq_4:address
	signal mm_interconnect_0_freq_3_s1_readdata                       : std_logic_vector(31 downto 0); -- freq_3:readdata -> mm_interconnect_0:freq_3_s1_readdata
	signal mm_interconnect_0_freq_3_s1_address                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:freq_3_s1_address -> freq_3:address
	signal mm_interconnect_0_freq_2_s1_readdata                       : std_logic_vector(31 downto 0); -- freq_2:readdata -> mm_interconnect_0:freq_2_s1_readdata
	signal mm_interconnect_0_freq_2_s1_address                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:freq_2_s1_address -> freq_2:address
	signal mm_interconnect_0_freq_1_s1_readdata                       : std_logic_vector(31 downto 0); -- freq_1:readdata -> mm_interconnect_0:freq_1_s1_readdata
	signal mm_interconnect_0_freq_1_s1_address                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:freq_1_s1_address -> freq_1:address
	signal mm_interconnect_0_freq_0_s1_readdata                       : std_logic_vector(31 downto 0); -- freq_0:readdata -> mm_interconnect_0:freq_0_s1_readdata
	signal mm_interconnect_0_freq_0_s1_address                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:freq_0_s1_address -> freq_0:address
	signal mm_interconnect_0_pwm_7_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:pwm_7_s1_chipselect -> pwm_7:chipselect
	signal mm_interconnect_0_pwm_7_s1_readdata                        : std_logic_vector(31 downto 0); -- pwm_7:readdata -> mm_interconnect_0:pwm_7_s1_readdata
	signal mm_interconnect_0_pwm_7_s1_address                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pwm_7_s1_address -> pwm_7:address
	signal mm_interconnect_0_pwm_7_s1_write                           : std_logic;                     -- mm_interconnect_0:pwm_7_s1_write -> mm_interconnect_0_pwm_7_s1_write:in
	signal mm_interconnect_0_pwm_7_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:pwm_7_s1_writedata -> pwm_7:writedata
	signal mm_interconnect_0_pwm_5_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:pwm_5_s1_chipselect -> pwm_5:chipselect
	signal mm_interconnect_0_pwm_5_s1_readdata                        : std_logic_vector(31 downto 0); -- pwm_5:readdata -> mm_interconnect_0:pwm_5_s1_readdata
	signal mm_interconnect_0_pwm_5_s1_address                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pwm_5_s1_address -> pwm_5:address
	signal mm_interconnect_0_pwm_5_s1_write                           : std_logic;                     -- mm_interconnect_0:pwm_5_s1_write -> mm_interconnect_0_pwm_5_s1_write:in
	signal mm_interconnect_0_pwm_5_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:pwm_5_s1_writedata -> pwm_5:writedata
	signal mm_interconnect_0_pwm_6_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:pwm_6_s1_chipselect -> pwm_6:chipselect
	signal mm_interconnect_0_pwm_6_s1_readdata                        : std_logic_vector(31 downto 0); -- pwm_6:readdata -> mm_interconnect_0:pwm_6_s1_readdata
	signal mm_interconnect_0_pwm_6_s1_address                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pwm_6_s1_address -> pwm_6:address
	signal mm_interconnect_0_pwm_6_s1_write                           : std_logic;                     -- mm_interconnect_0:pwm_6_s1_write -> mm_interconnect_0_pwm_6_s1_write:in
	signal mm_interconnect_0_pwm_6_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:pwm_6_s1_writedata -> pwm_6:writedata
	signal mm_interconnect_0_pwm_4_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:pwm_4_s1_chipselect -> pwm_4:chipselect
	signal mm_interconnect_0_pwm_4_s1_readdata                        : std_logic_vector(31 downto 0); -- pwm_4:readdata -> mm_interconnect_0:pwm_4_s1_readdata
	signal mm_interconnect_0_pwm_4_s1_address                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pwm_4_s1_address -> pwm_4:address
	signal mm_interconnect_0_pwm_4_s1_write                           : std_logic;                     -- mm_interconnect_0:pwm_4_s1_write -> mm_interconnect_0_pwm_4_s1_write:in
	signal mm_interconnect_0_pwm_4_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:pwm_4_s1_writedata -> pwm_4:writedata
	signal mm_interconnect_0_pwm_3_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:pwm_3_s1_chipselect -> pwm_3:chipselect
	signal mm_interconnect_0_pwm_3_s1_readdata                        : std_logic_vector(31 downto 0); -- pwm_3:readdata -> mm_interconnect_0:pwm_3_s1_readdata
	signal mm_interconnect_0_pwm_3_s1_address                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pwm_3_s1_address -> pwm_3:address
	signal mm_interconnect_0_pwm_3_s1_write                           : std_logic;                     -- mm_interconnect_0:pwm_3_s1_write -> mm_interconnect_0_pwm_3_s1_write:in
	signal mm_interconnect_0_pwm_3_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:pwm_3_s1_writedata -> pwm_3:writedata
	signal mm_interconnect_0_pwm_2_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:pwm_2_s1_chipselect -> pwm_2:chipselect
	signal mm_interconnect_0_pwm_2_s1_readdata                        : std_logic_vector(31 downto 0); -- pwm_2:readdata -> mm_interconnect_0:pwm_2_s1_readdata
	signal mm_interconnect_0_pwm_2_s1_address                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pwm_2_s1_address -> pwm_2:address
	signal mm_interconnect_0_pwm_2_s1_write                           : std_logic;                     -- mm_interconnect_0:pwm_2_s1_write -> mm_interconnect_0_pwm_2_s1_write:in
	signal mm_interconnect_0_pwm_2_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:pwm_2_s1_writedata -> pwm_2:writedata
	signal mm_interconnect_0_pwm_1_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:pwm_1_s1_chipselect -> pwm_1:chipselect
	signal mm_interconnect_0_pwm_1_s1_readdata                        : std_logic_vector(31 downto 0); -- pwm_1:readdata -> mm_interconnect_0:pwm_1_s1_readdata
	signal mm_interconnect_0_pwm_1_s1_address                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pwm_1_s1_address -> pwm_1:address
	signal mm_interconnect_0_pwm_1_s1_write                           : std_logic;                     -- mm_interconnect_0:pwm_1_s1_write -> mm_interconnect_0_pwm_1_s1_write:in
	signal mm_interconnect_0_pwm_1_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:pwm_1_s1_writedata -> pwm_1:writedata
	signal mm_interconnect_0_pwm_0_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:pwm_0_s1_chipselect -> pwm_0:chipselect
	signal mm_interconnect_0_pwm_0_s1_readdata                        : std_logic_vector(31 downto 0); -- pwm_0:readdata -> mm_interconnect_0:pwm_0_s1_readdata
	signal mm_interconnect_0_pwm_0_s1_address                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pwm_0_s1_address -> pwm_0:address
	signal mm_interconnect_0_pwm_0_s1_write                           : std_logic;                     -- mm_interconnect_0:pwm_0_s1_write -> mm_interconnect_0_pwm_0_s1_write:in
	signal mm_interconnect_0_pwm_0_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:pwm_0_s1_writedata -> pwm_0:writedata
	signal mm_interconnect_0_uart_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:uart_s1_chipselect -> uart:chipselect
	signal mm_interconnect_0_uart_s1_readdata                         : std_logic_vector(15 downto 0); -- uart:readdata -> mm_interconnect_0:uart_s1_readdata
	signal mm_interconnect_0_uart_s1_address                          : std_logic_vector(2 downto 0);  -- mm_interconnect_0:uart_s1_address -> uart:address
	signal mm_interconnect_0_uart_s1_read                             : std_logic;                     -- mm_interconnect_0:uart_s1_read -> mm_interconnect_0_uart_s1_read:in
	signal mm_interconnect_0_uart_s1_begintransfer                    : std_logic;                     -- mm_interconnect_0:uart_s1_begintransfer -> uart:begintransfer
	signal mm_interconnect_0_uart_s1_write                            : std_logic;                     -- mm_interconnect_0:uart_s1_write -> mm_interconnect_0_uart_s1_write:in
	signal mm_interconnect_0_uart_s1_writedata                        : std_logic_vector(15 downto 0); -- mm_interconnect_0:uart_s1_writedata -> uart:writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_chipselect           : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	signal mm_interconnect_0_onchip_memory2_0_s1_readdata             : std_logic_vector(31 downto 0); -- onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	signal mm_interconnect_0_onchip_memory2_0_s1_address              : std_logic_vector(11 downto 0); -- mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	signal mm_interconnect_0_onchip_memory2_0_s1_byteenable           : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	signal mm_interconnect_0_onchip_memory2_0_s1_write                : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	signal mm_interconnect_0_onchip_memory2_0_s1_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_clken                : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	signal mm_interconnect_0_tem_s1_readdata                          : std_logic_vector(31 downto 0); -- Tem:readdata -> mm_interconnect_0:Tem_s1_readdata
	signal mm_interconnect_0_tem_s1_address                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:Tem_s1_address -> Tem:address
	signal mm_interconnect_0_hum_s1_readdata                          : std_logic_vector(31 downto 0); -- Hum:readdata -> mm_interconnect_0:Hum_s1_readdata
	signal mm_interconnect_0_hum_s1_address                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:Hum_s1_address -> Hum:address
	signal irq_mapper_receiver0_irq                                   : std_logic;                     -- uart:irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                   : std_logic;                     -- timer_0:irq -> irq_mapper:receiver1_irq
	signal nios2_gen2_0_irq_irq                                       : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_gen2_0:irq
	signal rst_controller_reset_out_reset                             : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                         : std_logic;                     -- rst_controller:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	signal mm_interconnect_0_timer_0_s1_write_ports_inv               : std_logic;                     -- mm_interconnect_0_timer_0_s1_write:inv -> timer_0:write_n
	signal mm_interconnect_0_pwm_7_s1_write_ports_inv                 : std_logic;                     -- mm_interconnect_0_pwm_7_s1_write:inv -> pwm_7:write_n
	signal mm_interconnect_0_pwm_5_s1_write_ports_inv                 : std_logic;                     -- mm_interconnect_0_pwm_5_s1_write:inv -> pwm_5:write_n
	signal mm_interconnect_0_pwm_6_s1_write_ports_inv                 : std_logic;                     -- mm_interconnect_0_pwm_6_s1_write:inv -> pwm_6:write_n
	signal mm_interconnect_0_pwm_4_s1_write_ports_inv                 : std_logic;                     -- mm_interconnect_0_pwm_4_s1_write:inv -> pwm_4:write_n
	signal mm_interconnect_0_pwm_3_s1_write_ports_inv                 : std_logic;                     -- mm_interconnect_0_pwm_3_s1_write:inv -> pwm_3:write_n
	signal mm_interconnect_0_pwm_2_s1_write_ports_inv                 : std_logic;                     -- mm_interconnect_0_pwm_2_s1_write:inv -> pwm_2:write_n
	signal mm_interconnect_0_pwm_1_s1_write_ports_inv                 : std_logic;                     -- mm_interconnect_0_pwm_1_s1_write:inv -> pwm_1:write_n
	signal mm_interconnect_0_pwm_0_s1_write_ports_inv                 : std_logic;                     -- mm_interconnect_0_pwm_0_s1_write:inv -> pwm_0:write_n
	signal mm_interconnect_0_uart_s1_read_ports_inv                   : std_logic;                     -- mm_interconnect_0_uart_s1_read:inv -> uart:read_n
	signal mm_interconnect_0_uart_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_0_uart_s1_write:inv -> uart:write_n
	signal rst_controller_reset_out_reset_ports_inv                   : std_logic;                     -- rst_controller_reset_out_reset:inv -> [Hum:reset_n, Tem:reset_n, freq_0:reset_n, freq_1:reset_n, freq_2:reset_n, freq_3:reset_n, freq_4:reset_n, freq_5:reset_n, freq_6:reset_n, freq_7:reset_n, nios2_gen2_0:reset_n, pwm_0:reset_n, pwm_1:reset_n, pwm_2:reset_n, pwm_3:reset_n, pwm_4:reset_n, pwm_5:reset_n, pwm_6:reset_n, pwm_7:reset_n, timer_0:reset_n, uart:reset_n]

begin

	hum : component core_Hum
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_hum_s1_address,         --                  s1.address
			readdata => mm_interconnect_0_hum_s1_readdata,        --                    .readdata
			in_port  => hum_export                                -- external_connection.export
		);

	tem : component core_Hum
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_tem_s1_address,         --                  s1.address
			readdata => mm_interconnect_0_tem_s1_readdata,        --                    .readdata
			in_port  => tem_export                                -- external_connection.export
		);

	freq_0 : component core_freq_0
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_freq_0_s1_address,      --                  s1.address
			readdata => mm_interconnect_0_freq_0_s1_readdata,     --                    .readdata
			in_port  => freq_0_external_connection_export         -- external_connection.export
		);

	freq_1 : component core_freq_0
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_freq_1_s1_address,      --                  s1.address
			readdata => mm_interconnect_0_freq_1_s1_readdata,     --                    .readdata
			in_port  => freq_1_external_connection_export         -- external_connection.export
		);

	freq_2 : component core_freq_0
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_freq_2_s1_address,      --                  s1.address
			readdata => mm_interconnect_0_freq_2_s1_readdata,     --                    .readdata
			in_port  => freq_2_external_connection_export         -- external_connection.export
		);

	freq_3 : component core_freq_0
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_freq_3_s1_address,      --                  s1.address
			readdata => mm_interconnect_0_freq_3_s1_readdata,     --                    .readdata
			in_port  => freq_3_external_connection_export         -- external_connection.export
		);

	freq_4 : component core_freq_0
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_freq_4_s1_address,      --                  s1.address
			readdata => mm_interconnect_0_freq_4_s1_readdata,     --                    .readdata
			in_port  => freq_4_external_connection_export         -- external_connection.export
		);

	freq_5 : component core_freq_0
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_freq_5_s1_address,      --                  s1.address
			readdata => mm_interconnect_0_freq_5_s1_readdata,     --                    .readdata
			in_port  => freq_5_external_connection_export         -- external_connection.export
		);

	freq_6 : component core_freq_0
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_freq_6_s1_address,      --                  s1.address
			readdata => mm_interconnect_0_freq_6_s1_readdata,     --                    .readdata
			in_port  => freq_6_external_connection_export         -- external_connection.export
		);

	freq_7 : component core_freq_0
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_freq_7_s1_address,      --                  s1.address
			readdata => mm_interconnect_0_freq_7_s1_readdata,     --                    .readdata
			in_port  => freq_7_external_connection_export         -- external_connection.export
		);

	nios2_gen2_0 : component core_nios2_gen2_0
		port map (
			clk                                 => clk_clk,                                                    --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,                   --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                         --                          .reset_req
			d_address                           => nios2_gen2_0_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_gen2_0_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_gen2_0_data_master_read,                              --                          .read
			d_readdata                          => nios2_gen2_0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_gen2_0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_gen2_0_data_master_write,                             --                          .write
			d_writedata                         => nios2_gen2_0_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios2_gen2_0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_gen2_0_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_gen2_0_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_gen2_0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_gen2_0_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => nios2_gen2_0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2_gen2_0_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                        -- custom_instruction_master.readra
		);

	onchip_memory2_0 : component core_onchip_memory2_0
		port map (
			clk        => clk_clk,                                          --   clk1.clk
			address    => mm_interconnect_0_onchip_memory2_0_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory2_0_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory2_0_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory2_0_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory2_0_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory2_0_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory2_0_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                   -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,               --       .reset_req
			freeze     => '0'                                               -- (terminated)
		);

	pwm_0 : component core_pwm_0
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_pwm_0_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pwm_0_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pwm_0_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pwm_0_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pwm_0_s1_readdata,        --                    .readdata
			out_port   => pwm_0_external_connection_export            -- external_connection.export
		);

	pwm_1 : component core_pwm_0
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_pwm_1_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pwm_1_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pwm_1_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pwm_1_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pwm_1_s1_readdata,        --                    .readdata
			out_port   => pwm_1_external_connection_export            -- external_connection.export
		);

	pwm_2 : component core_pwm_0
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_pwm_2_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pwm_2_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pwm_2_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pwm_2_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pwm_2_s1_readdata,        --                    .readdata
			out_port   => pwm_2_external_connection_export            -- external_connection.export
		);

	pwm_3 : component core_pwm_0
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_pwm_3_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pwm_3_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pwm_3_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pwm_3_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pwm_3_s1_readdata,        --                    .readdata
			out_port   => pwm_3_external_connection_export            -- external_connection.export
		);

	pwm_4 : component core_pwm_0
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_pwm_4_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pwm_4_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pwm_4_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pwm_4_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pwm_4_s1_readdata,        --                    .readdata
			out_port   => pwm_4_external_connection_export            -- external_connection.export
		);

	pwm_5 : component core_pwm_0
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_pwm_5_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pwm_5_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pwm_5_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pwm_5_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pwm_5_s1_readdata,        --                    .readdata
			out_port   => pwm_5_external_connection_export            -- external_connection.export
		);

	pwm_6 : component core_pwm_0
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_pwm_6_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pwm_6_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pwm_6_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pwm_6_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pwm_6_s1_readdata,        --                    .readdata
			out_port   => pwm_6_external_connection_export            -- external_connection.export
		);

	pwm_7 : component core_pwm_0
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_pwm_7_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pwm_7_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pwm_7_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pwm_7_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pwm_7_s1_readdata,        --                    .readdata
			out_port   => pwm_7_external_connection_export            -- external_connection.export
		);

	timer_0 : component core_timer_0
		port map (
			clk        => clk_clk,                                      --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     -- reset.reset_n
			address    => mm_interconnect_0_timer_0_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_0_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_0_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_0_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_0_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver1_irq                      --   irq.irq
		);

	uart : component core_uart
		port map (
			clk           => clk_clk,                                   --                 clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address       => mm_interconnect_0_uart_s1_address,         --                  s1.address
			begintransfer => mm_interconnect_0_uart_s1_begintransfer,   --                    .begintransfer
			chipselect    => mm_interconnect_0_uart_s1_chipselect,      --                    .chipselect
			read_n        => mm_interconnect_0_uart_s1_read_ports_inv,  --                    .read_n
			write_n       => mm_interconnect_0_uart_s1_write_ports_inv, --                    .write_n
			writedata     => mm_interconnect_0_uart_s1_writedata,       --                    .writedata
			readdata      => mm_interconnect_0_uart_s1_readdata,        --                    .readdata
			rxd           => uart_external_connection_rxd,              -- external_connection.export
			txd           => uart_external_connection_txd,              --                    .export
			irq           => irq_mapper_receiver0_irq                   --                 irq.irq
		);

	mm_interconnect_0 : component core_mm_interconnect_0
		port map (
			clk_0_clk_clk                                  => clk_clk,                                                    --                                clk_0_clk.clk
			nios2_gen2_0_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                             -- nios2_gen2_0_reset_reset_bridge_in_reset.reset
			nios2_gen2_0_data_master_address               => nios2_gen2_0_data_master_address,                           --                 nios2_gen2_0_data_master.address
			nios2_gen2_0_data_master_waitrequest           => nios2_gen2_0_data_master_waitrequest,                       --                                         .waitrequest
			nios2_gen2_0_data_master_byteenable            => nios2_gen2_0_data_master_byteenable,                        --                                         .byteenable
			nios2_gen2_0_data_master_read                  => nios2_gen2_0_data_master_read,                              --                                         .read
			nios2_gen2_0_data_master_readdata              => nios2_gen2_0_data_master_readdata,                          --                                         .readdata
			nios2_gen2_0_data_master_write                 => nios2_gen2_0_data_master_write,                             --                                         .write
			nios2_gen2_0_data_master_writedata             => nios2_gen2_0_data_master_writedata,                         --                                         .writedata
			nios2_gen2_0_data_master_debugaccess           => nios2_gen2_0_data_master_debugaccess,                       --                                         .debugaccess
			nios2_gen2_0_instruction_master_address        => nios2_gen2_0_instruction_master_address,                    --          nios2_gen2_0_instruction_master.address
			nios2_gen2_0_instruction_master_waitrequest    => nios2_gen2_0_instruction_master_waitrequest,                --                                         .waitrequest
			nios2_gen2_0_instruction_master_read           => nios2_gen2_0_instruction_master_read,                       --                                         .read
			nios2_gen2_0_instruction_master_readdata       => nios2_gen2_0_instruction_master_readdata,                   --                                         .readdata
			freq_0_s1_address                              => mm_interconnect_0_freq_0_s1_address,                        --                                freq_0_s1.address
			freq_0_s1_readdata                             => mm_interconnect_0_freq_0_s1_readdata,                       --                                         .readdata
			freq_1_s1_address                              => mm_interconnect_0_freq_1_s1_address,                        --                                freq_1_s1.address
			freq_1_s1_readdata                             => mm_interconnect_0_freq_1_s1_readdata,                       --                                         .readdata
			freq_2_s1_address                              => mm_interconnect_0_freq_2_s1_address,                        --                                freq_2_s1.address
			freq_2_s1_readdata                             => mm_interconnect_0_freq_2_s1_readdata,                       --                                         .readdata
			freq_3_s1_address                              => mm_interconnect_0_freq_3_s1_address,                        --                                freq_3_s1.address
			freq_3_s1_readdata                             => mm_interconnect_0_freq_3_s1_readdata,                       --                                         .readdata
			freq_4_s1_address                              => mm_interconnect_0_freq_4_s1_address,                        --                                freq_4_s1.address
			freq_4_s1_readdata                             => mm_interconnect_0_freq_4_s1_readdata,                       --                                         .readdata
			freq_5_s1_address                              => mm_interconnect_0_freq_5_s1_address,                        --                                freq_5_s1.address
			freq_5_s1_readdata                             => mm_interconnect_0_freq_5_s1_readdata,                       --                                         .readdata
			freq_6_s1_address                              => mm_interconnect_0_freq_6_s1_address,                        --                                freq_6_s1.address
			freq_6_s1_readdata                             => mm_interconnect_0_freq_6_s1_readdata,                       --                                         .readdata
			freq_7_s1_address                              => mm_interconnect_0_freq_7_s1_address,                        --                                freq_7_s1.address
			freq_7_s1_readdata                             => mm_interconnect_0_freq_7_s1_readdata,                       --                                         .readdata
			Hum_s1_address                                 => mm_interconnect_0_hum_s1_address,                           --                                   Hum_s1.address
			Hum_s1_readdata                                => mm_interconnect_0_hum_s1_readdata,                          --                                         .readdata
			nios2_gen2_0_debug_mem_slave_address           => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,     --             nios2_gen2_0_debug_mem_slave.address
			nios2_gen2_0_debug_mem_slave_write             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,       --                                         .write
			nios2_gen2_0_debug_mem_slave_read              => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,        --                                         .read
			nios2_gen2_0_debug_mem_slave_readdata          => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,    --                                         .readdata
			nios2_gen2_0_debug_mem_slave_writedata         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,   --                                         .writedata
			nios2_gen2_0_debug_mem_slave_byteenable        => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,  --                                         .byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest       => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest, --                                         .waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess       => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess, --                                         .debugaccess
			onchip_memory2_0_s1_address                    => mm_interconnect_0_onchip_memory2_0_s1_address,              --                      onchip_memory2_0_s1.address
			onchip_memory2_0_s1_write                      => mm_interconnect_0_onchip_memory2_0_s1_write,                --                                         .write
			onchip_memory2_0_s1_readdata                   => mm_interconnect_0_onchip_memory2_0_s1_readdata,             --                                         .readdata
			onchip_memory2_0_s1_writedata                  => mm_interconnect_0_onchip_memory2_0_s1_writedata,            --                                         .writedata
			onchip_memory2_0_s1_byteenable                 => mm_interconnect_0_onchip_memory2_0_s1_byteenable,           --                                         .byteenable
			onchip_memory2_0_s1_chipselect                 => mm_interconnect_0_onchip_memory2_0_s1_chipselect,           --                                         .chipselect
			onchip_memory2_0_s1_clken                      => mm_interconnect_0_onchip_memory2_0_s1_clken,                --                                         .clken
			pwm_0_s1_address                               => mm_interconnect_0_pwm_0_s1_address,                         --                                 pwm_0_s1.address
			pwm_0_s1_write                                 => mm_interconnect_0_pwm_0_s1_write,                           --                                         .write
			pwm_0_s1_readdata                              => mm_interconnect_0_pwm_0_s1_readdata,                        --                                         .readdata
			pwm_0_s1_writedata                             => mm_interconnect_0_pwm_0_s1_writedata,                       --                                         .writedata
			pwm_0_s1_chipselect                            => mm_interconnect_0_pwm_0_s1_chipselect,                      --                                         .chipselect
			pwm_1_s1_address                               => mm_interconnect_0_pwm_1_s1_address,                         --                                 pwm_1_s1.address
			pwm_1_s1_write                                 => mm_interconnect_0_pwm_1_s1_write,                           --                                         .write
			pwm_1_s1_readdata                              => mm_interconnect_0_pwm_1_s1_readdata,                        --                                         .readdata
			pwm_1_s1_writedata                             => mm_interconnect_0_pwm_1_s1_writedata,                       --                                         .writedata
			pwm_1_s1_chipselect                            => mm_interconnect_0_pwm_1_s1_chipselect,                      --                                         .chipselect
			pwm_2_s1_address                               => mm_interconnect_0_pwm_2_s1_address,                         --                                 pwm_2_s1.address
			pwm_2_s1_write                                 => mm_interconnect_0_pwm_2_s1_write,                           --                                         .write
			pwm_2_s1_readdata                              => mm_interconnect_0_pwm_2_s1_readdata,                        --                                         .readdata
			pwm_2_s1_writedata                             => mm_interconnect_0_pwm_2_s1_writedata,                       --                                         .writedata
			pwm_2_s1_chipselect                            => mm_interconnect_0_pwm_2_s1_chipselect,                      --                                         .chipselect
			pwm_3_s1_address                               => mm_interconnect_0_pwm_3_s1_address,                         --                                 pwm_3_s1.address
			pwm_3_s1_write                                 => mm_interconnect_0_pwm_3_s1_write,                           --                                         .write
			pwm_3_s1_readdata                              => mm_interconnect_0_pwm_3_s1_readdata,                        --                                         .readdata
			pwm_3_s1_writedata                             => mm_interconnect_0_pwm_3_s1_writedata,                       --                                         .writedata
			pwm_3_s1_chipselect                            => mm_interconnect_0_pwm_3_s1_chipselect,                      --                                         .chipselect
			pwm_4_s1_address                               => mm_interconnect_0_pwm_4_s1_address,                         --                                 pwm_4_s1.address
			pwm_4_s1_write                                 => mm_interconnect_0_pwm_4_s1_write,                           --                                         .write
			pwm_4_s1_readdata                              => mm_interconnect_0_pwm_4_s1_readdata,                        --                                         .readdata
			pwm_4_s1_writedata                             => mm_interconnect_0_pwm_4_s1_writedata,                       --                                         .writedata
			pwm_4_s1_chipselect                            => mm_interconnect_0_pwm_4_s1_chipselect,                      --                                         .chipselect
			pwm_5_s1_address                               => mm_interconnect_0_pwm_5_s1_address,                         --                                 pwm_5_s1.address
			pwm_5_s1_write                                 => mm_interconnect_0_pwm_5_s1_write,                           --                                         .write
			pwm_5_s1_readdata                              => mm_interconnect_0_pwm_5_s1_readdata,                        --                                         .readdata
			pwm_5_s1_writedata                             => mm_interconnect_0_pwm_5_s1_writedata,                       --                                         .writedata
			pwm_5_s1_chipselect                            => mm_interconnect_0_pwm_5_s1_chipselect,                      --                                         .chipselect
			pwm_6_s1_address                               => mm_interconnect_0_pwm_6_s1_address,                         --                                 pwm_6_s1.address
			pwm_6_s1_write                                 => mm_interconnect_0_pwm_6_s1_write,                           --                                         .write
			pwm_6_s1_readdata                              => mm_interconnect_0_pwm_6_s1_readdata,                        --                                         .readdata
			pwm_6_s1_writedata                             => mm_interconnect_0_pwm_6_s1_writedata,                       --                                         .writedata
			pwm_6_s1_chipselect                            => mm_interconnect_0_pwm_6_s1_chipselect,                      --                                         .chipselect
			pwm_7_s1_address                               => mm_interconnect_0_pwm_7_s1_address,                         --                                 pwm_7_s1.address
			pwm_7_s1_write                                 => mm_interconnect_0_pwm_7_s1_write,                           --                                         .write
			pwm_7_s1_readdata                              => mm_interconnect_0_pwm_7_s1_readdata,                        --                                         .readdata
			pwm_7_s1_writedata                             => mm_interconnect_0_pwm_7_s1_writedata,                       --                                         .writedata
			pwm_7_s1_chipselect                            => mm_interconnect_0_pwm_7_s1_chipselect,                      --                                         .chipselect
			Tem_s1_address                                 => mm_interconnect_0_tem_s1_address,                           --                                   Tem_s1.address
			Tem_s1_readdata                                => mm_interconnect_0_tem_s1_readdata,                          --                                         .readdata
			timer_0_s1_address                             => mm_interconnect_0_timer_0_s1_address,                       --                               timer_0_s1.address
			timer_0_s1_write                               => mm_interconnect_0_timer_0_s1_write,                         --                                         .write
			timer_0_s1_readdata                            => mm_interconnect_0_timer_0_s1_readdata,                      --                                         .readdata
			timer_0_s1_writedata                           => mm_interconnect_0_timer_0_s1_writedata,                     --                                         .writedata
			timer_0_s1_chipselect                          => mm_interconnect_0_timer_0_s1_chipselect,                    --                                         .chipselect
			uart_s1_address                                => mm_interconnect_0_uart_s1_address,                          --                                  uart_s1.address
			uart_s1_write                                  => mm_interconnect_0_uart_s1_write,                            --                                         .write
			uart_s1_read                                   => mm_interconnect_0_uart_s1_read,                             --                                         .read
			uart_s1_readdata                               => mm_interconnect_0_uart_s1_readdata,                         --                                         .readdata
			uart_s1_writedata                              => mm_interconnect_0_uart_s1_writedata,                        --                                         .writedata
			uart_s1_begintransfer                          => mm_interconnect_0_uart_s1_begintransfer,                    --                                         .begintransfer
			uart_s1_chipselect                             => mm_interconnect_0_uart_s1_chipselect                        --                                         .chipselect
		);

	irq_mapper : component core_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			sender_irq    => nios2_gen2_0_irq_irq            --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => nios2_gen2_0_debug_reset_request_reset, -- reset_in0.reset
			reset_in1      => nios2_gen2_0_debug_reset_request_reset, -- reset_in1.reset
			clk            => clk_clk,                                --       clk.clk
			reset_out      => rst_controller_reset_out_reset,         -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,     --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	mm_interconnect_0_timer_0_s1_write_ports_inv <= not mm_interconnect_0_timer_0_s1_write;

	mm_interconnect_0_pwm_7_s1_write_ports_inv <= not mm_interconnect_0_pwm_7_s1_write;

	mm_interconnect_0_pwm_5_s1_write_ports_inv <= not mm_interconnect_0_pwm_5_s1_write;

	mm_interconnect_0_pwm_6_s1_write_ports_inv <= not mm_interconnect_0_pwm_6_s1_write;

	mm_interconnect_0_pwm_4_s1_write_ports_inv <= not mm_interconnect_0_pwm_4_s1_write;

	mm_interconnect_0_pwm_3_s1_write_ports_inv <= not mm_interconnect_0_pwm_3_s1_write;

	mm_interconnect_0_pwm_2_s1_write_ports_inv <= not mm_interconnect_0_pwm_2_s1_write;

	mm_interconnect_0_pwm_1_s1_write_ports_inv <= not mm_interconnect_0_pwm_1_s1_write;

	mm_interconnect_0_pwm_0_s1_write_ports_inv <= not mm_interconnect_0_pwm_0_s1_write;

	mm_interconnect_0_uart_s1_read_ports_inv <= not mm_interconnect_0_uart_s1_read;

	mm_interconnect_0_uart_s1_write_ports_inv <= not mm_interconnect_0_uart_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of core
